/*
[TB_INFO_START]
Name: tb_uart_ascii_sender
Target: uart_ascii_sender
Role: Testbench for ASCII Report Generator
Scenario:
  - Stimulates request inputs for Watch, SR04, DHT11, and Loopback
  - Assumes TX FIFO is always ready (no full backpressure)
CheckPoint:
  - Captures serialized UART output into a log
  - Verifies correct formatting of strings (e.g., "WATCH...", "TEMP...")
  - Checks arbitration priority if multiple requests occur
[TB_INFO_END]
*/

`timescale 1ns / 1ps

module tb_uart_ascii_sender;
  // initial begin
  //   $dumpfile("tb_uart_ascii_sender.vcd");
  //   $dumpvars(0, tb_uart_ascii_sender);
  // end

  reg iClk;
  reg iRst;

  wire iTxFifoFull;
  wire [7:0] oTxData;
  wire oTxPushValid;

  reg [7:0] iLoopData;
  reg iLoopValid;
  reg iReqWatchReport;
  reg iReqSr04Report;
  reg iReqTempReport;
  reg iReqHumReport;
  reg [6:0] iWatchHour, iWatchMin, iWatchSec;
  reg [9:0] iSr04DistanceCm;
  reg iSr04DistanceValid;
  reg [7:0] iDhtHumInt;
  reg [7:0] iDhtTempInt;
  reg iDhtDataValid;

  uart_ascii_sender dut (
    .iClk(iClk),
    .iRst(iRst),
    .iTxFifoFull(iTxFifoFull),
    .oTxData(oTxData),
    .oTxPushValid(oTxPushValid),
    .iLoopData(iLoopData),
    .iLoopValid(iLoopValid),
    .iReqWatchReport(iReqWatchReport),
    .iReqSr04Report(iReqSr04Report),
    .iReqTempReport(iReqTempReport),
    .iReqHumReport(iReqHumReport),
    .iWatchHour(iWatchHour),
    .iWatchMin(iWatchMin),
    .iWatchSec(iWatchSec),
    .iSr04DistanceCm(iSr04DistanceCm),
    .iSr04DistanceValid(iSr04DistanceValid),
    .iDhtHumInt(iDhtHumInt),
    .iDhtTempInt(iDhtTempInt),
    .iDhtDataValid(iDhtDataValid)
  );

  always #5 iClk = ~iClk;
  assign iTxFifoFull = 1'b0;

  integer i;
  reg [7:0] tx_count;
  reg [7:0] tx_log [0:255];
  // Expected bytes for this stimulus:
  // 1(loop) + 18(watch) + 14(sr04) + 12(temp) + 11(hum) = 56
  localparam [7:0] EXP_TX_COUNT = 8'd56;

  always @(posedge iClk or posedge iRst) begin
    if (iRst) begin
      tx_count <= 8'h0;
      for(i=0;i<256;i=i+1) begin
        tx_log[i] <= 8'h0;
      end 
    end 
    else begin
      if (oTxPushValid) begin
        tx_log[tx_count] <= oTxData;
        tx_count <= tx_count + 8'd1;
      end
    end
  end

  task pulse_loop(input [7:0] ch);
    begin
      @(posedge iClk);
      iLoopData  <= ch;
      iLoopValid <= 1'b1;
      @(posedge iClk);
      iLoopValid <= 1'b0;
    end
  endtask

  task pulse_watch_report;
    begin
      @(posedge iClk);
      iReqWatchReport <= 1'b1;
      @(posedge iClk);
      iReqWatchReport <= 1'b0;
    end
  endtask

  task pulse_sr04_report;
    begin
      @(posedge iClk);
      iReqSr04Report <= 1'b1;
      @(posedge iClk);
      iReqSr04Report <= 1'b0;
    end
  endtask

  task pulse_temp_report;
    begin
      @(posedge iClk);
      iReqTempReport <= 1'b1;
      @(posedge iClk);
      iReqTempReport <= 1'b0;
    end
  endtask

  task pulse_hum_report;
    begin
      @(posedge iClk);
      iReqHumReport <= 1'b1;
      @(posedge iClk);
      iReqHumReport <= 1'b0;
    end
  endtask

  initial begin
    iClk = 1'b0;
    iRst = 1'b1;

    iLoopData = 8'd0;
    iLoopValid = 1'b0;
    iReqWatchReport = 1'b0;
    iReqSr04Report = 1'b0;
    iReqTempReport = 1'b0;
    iReqHumReport = 1'b0;

    iWatchHour = 7'd12;
    iWatchMin  = 7'd34;
    iWatchSec  = 7'd56;
    iSr04DistanceCm = 10'd123;
    iSr04DistanceValid = 1'b1;
    iDhtHumInt = 8'd44;
    iDhtTempInt = 8'd23;
    iDhtDataValid = 1'b1;

    repeat (5) @(posedge iClk);
    iRst = 1'b0;

    pulse_loop("A");//loopback test
    pulse_watch_report();
    pulse_sr04_report();
    pulse_temp_report();
    pulse_hum_report();

    wait (tx_count == EXP_TX_COUNT);
    repeat (10) @(posedge iClk);
    // // Extra guard: ensure no unexpected additional bytes.
    // 
    // if (tx_count !== EXP_TX_COUNT) begin
    //   $display("uart_ascii_sender extra bytes detected: exp=%0d act=%0d", EXP_TX_COUNT, tx_count);
    //   $finish;
    // end

    $display("tb_uart_ascii_sender finished: tx_count=%0d", tx_count);
    for (i = 0; i < tx_count; i = i + 1) begin
      if (tx_log[i] == 8'h0D) begin
        $display("tx_log[%0d] = 0x%02h (CR)", i, tx_log[i]);
      end else if (tx_log[i] == 8'h0A) begin
        $display("tx_log[%0d] = 0x%02h (LF)", i, tx_log[i]);
      end else if ((tx_log[i] >= 8'h20) && (tx_log[i] <= 8'h7E)) begin
        $display("tx_log[%0d] = 0x%02h (%c)", i, tx_log[i], tx_log[i]);
      end else begin
        $display("tx_log[%0d] = 0x%02h (.)", i, tx_log[i]);
      end
    end
    $finish;
  end

endmodule
